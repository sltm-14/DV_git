
`ifndef ROOT_SV
    `define ROOT_SV
module root
import system_mdr_pkg::*;
(
	input clk,
	input reset,
	input i_enable,
	input i_dataX,
	
	output data_t o_quotation,
	output data_t o_remainder
);


	

endmodule
`endif