library verilog;
use verilog.vl_types.all;
entity clk_pkg is
end clk_pkg;
