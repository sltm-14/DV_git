library verilog;
use verilog.vl_types.all;
entity switch_pkg is
end switch_pkg;
