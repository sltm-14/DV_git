library verilog;
use verilog.vl_types.all;
entity compA2_data is
end compA2_data;
