library verilog;
use verilog.vl_types.all;
entity tb_siso_left is
end tb_siso_left;
