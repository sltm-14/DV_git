`ifndef MUX_DATA_SV
    `define MUX_DATA_SV

module mux_data
import pkg_system_mdr::*;(
	if_mdr.mux_data mux
	);

	

endmodule