`ifndef SYSTEM_MDR_PKG_SV
    `define SYSTEM_MDR_PKG_SV
package system_mdr_pkg;

    localparam  DW      	= 16;

    typedef logic [DW-1:0]		data_t;
    typedef logic [1:0]			enb_t;

endpackage

`endif
