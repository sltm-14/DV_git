library verilog;
use verilog.vl_types.all;
entity add_con is
    port(
        i_hto_0         : in     vl_logic;
        i_hto_1         : in     vl_logic;
        i_hto_2         : in     vl_logic;
        i_hto_3         : in     vl_logic;
        o_hto_0         : out    vl_logic;
        o_hto_1         : out    vl_logic;
        o_hto_2         : out    vl_logic;
        o_hto_3         : out    vl_logic
    );
end add_con;
