library verilog;
use verilog.vl_types.all;
entity pkg_mult is
end pkg_mult;
