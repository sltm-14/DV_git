`ifndef QUOTIENT_SV
    `define QUOTIENT_SV

module quotient
import pkg_system_mdr::*;(

	);

endmodule