library verilog;
use verilog.vl_types.all;
entity leds_pkg is
end leds_pkg;
