`ifndef CONTROL_SV
    `define CONTROL_SV

module control
import mxv_pkg::*;
(
	input clk_wr,
	input clk_rd,
	input rst,

	input data_uart_t data,


);

endmodule
`endif