`ifndef MUX_REMINDER_SV
    `define MUX_REMINDER_SV

module mux_reminder
import pkg_system_mdr::*;(

	);

endmodule