`ifndef REMINDER_SV
    `define REMINDER_SV

module reminder
import pkg_system_mdr::*;(

	);

endmodule