`ifndef MUX_OR_SV
    `define MUX_OR_SV

module mux_or
import pkg_system_mdr::*;(

	);

endmodule