library verilog;
use verilog.vl_types.all;
entity tb_ms is
end tb_ms;
