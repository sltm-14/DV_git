library verilog;
use verilog.vl_types.all;
entity pkg_bin_to_thto is
end pkg_bin_to_thto;
