library verilog;
use verilog.vl_types.all;
entity mult_pkg is
end mult_pkg;
