library verilog;
use verilog.vl_types.all;
entity comp2_pkg is
end comp2_pkg;
