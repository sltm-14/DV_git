`ifndef MUX_QUOTIENT_SV
    `define MUX_QUOTIENT_SV

module mux_quotinet
import pkg_system_mdr::*;(

	);

endmodule