/*-----------------------------------------------
* MODULE: 	  	display_if.sv
* DESCRIPTION: Interface with modports of the
*					display the modules					
*					error
* VERSION:    	1.0
* AUTHORS:    	Andres Hernandez, Carem Acosta
* DATE:       	05 / 04 / 19
* ----------------------------------------------*/
`ifndef DISPLAY_IF_SV
	`define DISPLAY_IF_SV

interface display_if();
import system_mdr_pkg::*;




endinterface

`endif