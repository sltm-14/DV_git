library verilog;
use verilog.vl_types.all;
entity ms is
    port(
        i_clk           : in     vl_logic;
        i_rst           : in     vl_logic;
        i_start         : in     vl_logic;
        i_sw0           : in     vl_logic;
        i_sw1           : in     vl_logic;
        i_sw2           : in     vl_logic;
        i_sw3           : in     vl_logic;
        i_sw4           : in     vl_logic;
        i_sw5           : in     vl_logic;
        i_sw6           : in     vl_logic;
        i_sw7           : in     vl_logic;
        i_sw8           : in     vl_logic;
        i_sw9           : in     vl_logic;
        i_sw10          : in     vl_logic;
        i_sw11          : in     vl_logic;
        i_sw12          : in     vl_logic;
        i_sw13          : in     vl_logic;
        i_sw14          : in     vl_logic;
        i_sw15          : in     vl_logic;
        i_sw16          : in     vl_logic;
        i_sw17          : in     vl_logic;
        o_led0          : out    vl_logic;
        o_led1          : out    vl_logic;
        o_led2          : out    vl_logic;
        o_led3          : out    vl_logic;
        o_led4          : out    vl_logic;
        o_led5          : out    vl_logic;
        o_led6          : out    vl_logic;
        o_led7          : out    vl_logic;
        o_led8          : out    vl_logic;
        o_led9          : out    vl_logic;
        o_led10         : out    vl_logic;
        o_led11         : out    vl_logic;
        o_led12         : out    vl_logic;
        o_led13         : out    vl_logic;
        o_led14         : out    vl_logic;
        o_led15         : out    vl_logic;
        o_led16         : out    vl_logic;
        o_ready         : out    vl_logic;
        test            : out    vl_logic
    );
end ms;
