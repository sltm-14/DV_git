library verilog;
use verilog.vl_types.all;
entity control_pkg is
end control_pkg;
