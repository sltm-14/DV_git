`ifndef COMPA2_DATA_SV
    `define COMPA2_DATA_SV

module compA2_data
import pkg_system_mdr::*;(

	);

endmodule 