library verilog;
use verilog.vl_types.all;
entity tb_piso_msb is
end tb_piso_msb;
