`ifndef MUX_B_SV
    `define MUX_B_SV

module mux_b
import pkg_system_mdr::*;(

	);

endmodule