library verilog;
use verilog.vl_types.all;
entity tb_sipo is
end tb_sipo;
