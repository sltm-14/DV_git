`ifndef MUX_A_SV
    `define MUX_A_SV

module mux_a
import pkg_system_mdr::*;(

	);

endmodule