`ifndef ALU_SV
    `define ALU_SV

module alu
import pkg_system_mdr::*;(

	);

endmodule 