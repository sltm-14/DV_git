library verilog;
use verilog.vl_types.all;
entity pkg_system_mdr is
end pkg_system_mdr;
