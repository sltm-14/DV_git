`ifndef COMPA2_QUOTIENT_SV
    `define COMPA2_QUOTIENT_SV

module compA2_quotient
import pkg_system_mdr::*;(

	);

endmodule 