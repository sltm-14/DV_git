`ifndef COMPA2_REMINDER_SV
    `define MDR_SV

module compA2_reminder
import pkg_system_mdr::*;(

	);

endmodule